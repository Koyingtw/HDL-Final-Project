module sender(clk, prefix, argc, argv1, argv2);
    input clk;
    input [7:0] prefix;
    input [7:0] argc;
    input [7:0] argv1;
    input [7:0] argv2;


    logic [7:0] queue [$:127];

    

endmodule